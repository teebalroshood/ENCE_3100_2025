module multiplier_8x8(
    input  [7:0]  i_A,
    input  [7:0]  i_B,
    output [15:0] o_P,
    output        o_Overflow
);
    // ----------------------------------------------------
    // Partial product generation (AND array)
    // ----------------------------------------------------
    wire [7:0] pp [7:0];
    genvar i;
    generate
        for (i = 0; i < 8; i = i + 1) begin : gen_pp
            assign pp[i] = i_A & {8{i_B[i]}};
        end
    endgenerate

    // ----------------------------------------------------
    // First Stage of Adders (add pp[0] and shifted pp[1])
    // ----------------------------------------------------
    wire [15:0] stage1 = {8'b0, pp[0]} + {7'b0, pp[1], 1'b0};

    // ----------------------------------------------------
    // Second Stage of Adders (add shifted pp[2])
    // ----------------------------------------------------
    wire [15:0] stage2 = stage1 + {6'b0, pp[2], 2'b0};

    // ----------------------------------------------------
    // Third Stage of Adders (add shifted pp[3])
    // ----------------------------------------------------
    wire [15:0] stage3 = stage2 + {5'b0, pp[3], 3'b0};

    // ----------------------------------------------------
    // Fourth Stage of Adders (add shifted pp[4])
    // ----------------------------------------------------
    wire [15:0] stage4 = stage3 + {4'b0, pp[4], 4'b0};

    // ----------------------------------------------------
    // Fifth Stage of Adders (add shifted pp[5])
    // ----------------------------------------------------
    wire [15:0] stage5 = stage4 + {3'b0, pp[5], 5'b0};

    // ----------------------------------------------------
    // Sixth Stage of Adders (add shifted pp[6])
    // ----------------------------------------------------
    wire [15:0] stage6 = stage5 + {2'b0, pp[6], 6'b0};

    // ----------------------------------------------------
    // Seventh Stage of Adders (add shifted pp[7])
    // ----------------------------------------------------
    wire [15:0] stage7 = stage6 + {1'b0, pp[7], 7'b0};

    // ----------------------------------------------------
    // Final Product
    // ----------------------------------------------------
    assign o_P = stage7;
    assign o_Overflow = |stage7[15:8];

endmodule
