module dff_posedge(input D, input Clk, input rst_n, output reg Q);
  always @(posedge Clk or negedge rst_n)
    if (!rst_n) Q <= 1'b0; else Q <= D;
endmodule