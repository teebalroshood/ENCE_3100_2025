// test.v

// Generated using ACDS version 24.1 1077

`timescale 1 ps / 1 ps
module test (
		input  wire [12:0] a,      //      a.a
		input  wire        areset, // areset.reset
		output wire [9:0]  c,      //      c.c
		input  wire        clk,    //    clk.clk
		input  wire [0:0]  en,     //     en.en
		output wire [9:0]  s       //      s.s
	);

	test_CORDIC_0 cordic_0 (
		.clk    (clk),    //    clk.clk
		.areset (areset), // areset.reset
		.en     (en),     //     en.en
		.a      (a),      //      a.a
		.c      (c),      //      c.c
		.s      (s)       //      s.s
	);

endmodule
